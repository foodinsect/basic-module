// Johnson Counter with Initial Value
// 2^N-2N invalid states and 2N valid states -> Half number of FF for same states
module johnson_counter #(
    parameter N = 4             // Define the default size of the counter
)(
    input wire clk,             // Clock signal
    input wire start,           // Start signal to initialize the counter
    output reg [0:N-1] qout     // Counter output
);
    

    // Counter logic
    always @(posedge clk or posedge start) begin
        if (start)
            qout <= {N{1'b0}};                  // Initialize counter with "0000"
        else
            qout <= {~qout[N-1], qout[0:N-2]};  // Shift left with inverted MSB at LSB
    end
endmodule
